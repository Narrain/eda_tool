module hello;
    logic a;
    logic b;
    assign b = a;
endmodule
