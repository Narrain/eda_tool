module top;
    wire a;
    assign a = 1'b1;
endmodule
